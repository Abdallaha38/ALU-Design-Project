LIBRARY iee;
USE iee.std_logic_1164.all;
